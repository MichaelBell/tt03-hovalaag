/* Copyright (C) 2023 Michael Bell

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
*/

/*
   Wrapper for the Hovalaag CPU.  This provides registers for the data coming in
   over the 6-bit in to populate, and exposes the outputs for the 8-bit output bus
   */

module HovalaagWrapper(
    input clk,     // Clock for the wrapper
    input reset_n,
    input reset_rosc_n,

    input [2:0] addr, // Input is DDR
                      // Input:  0-2: Set instr bits 0-5, 6-11, 12-17, 18-23, 24-29, 30-31
                      //           3: Set IN1 bits 0-5, 6-11  
                      //           4: Set IN2 bits 0-5, 6-11
                      // Output:   2: Execute status: 0: IN1 advance, 1: IN2 advance, 2: OUT1 valid, 3: OUT2 valid
                      //           4: New PC
                      //           0-1: OUT bits 0-7, 8-11 (valid for OUT1 or OUT2 if one of the valid bits was set)
                      //           3: OUT bits 0-3, 11 in 7-segment format (11 sets the 8th output)
    input [5:0] io_in,
    output [7:0] io_out
);
    reg [31:0] instr;
    reg [11:0] in1;
    reg [11:0] in2;

    wire in1_adv;
    wire in2_adv;
    wire [11:0] out;
    wire out_valid;
    wire out_select;
    wire [7:0] pc;

    wire [5:0] fast_count;
    reg [5:0] buffered_fast_count;
    reg [11:0] rng_bits;

    wire [6:0] seg7_out;

    Hovalaag hov (
        .clk(clk),
        .clk_en(addr == 3),
        .IN1(in1),
        .IN1_adv(in1_adv),
        .IN2(in2),
        .IN2_adv(in2_adv),
        .OUT(out),
        .instr(instr),
        .PC_out(pc),
        .rst(!reset_n),
        .alu_op_14_source(rng_bits),
        .alu_op_15_source(12'h001)
    );

    Seg7 seg7 (
        .value(out[3:0]),
        .seg_out(seg7_out)
    );

    reg rosc_pause;

    RingOscillator #(.NUM_FAST_CLKS(6), .STAGES(11)) rosc (
        .reset_n(reset_rosc_n),
        .pause(rosc_pause),
        .fast_clk(fast_count)
    );

    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            rosc_pause <= 1'b0;
            rng_bits <= 0;
        end else begin
            if (rosc_pause) begin
                rng_bits[11:6] <= rng_bits[5:0];
                rng_bits[5:0] <= buffered_fast_count[5:0];
            end
            rosc_pause <= ~rosc_pause;
        end
    end

`ifdef SIM
    always @(negedge clk) begin
        buffered_fast_count[5:0] <= fast_count & {6{rosc_pause}};
    end
`else
    genvar i;
    generate
        for (i = 0; i < 6; i = i + 1) begin
            sky130_fd_sc_hd__dlrtn_1 fastcntlatch(.Q(buffered_fast_count[i]), .D(fast_count[i] && rosc_pause), .GATE_N(clk), .RESET_B(reset_n));
        end
    endgenerate
`endif

    // We want to use out valid and select before the result is clocked out,
    // so decode them directly here
    assign out_valid = instr[14];
    assign out_select = instr[13];

    always @(posedge clk) begin
        if (!reset_n) begin
            instr[5:0] <= 0;
            instr[17:12] <= 0;
            instr[29:24] <= 0;
            in1[5:0] <= 0;
            in2[5:0] <= 0;
        end
        else begin
            case (addr)
            0: instr[ 5: 0] <= io_in;
            1: instr[17:12] <= io_in;
            2: instr[29:24] <= io_in;
            3: in1[5: 0] <= io_in;
            4: in2[5: 0] <= io_in;
            endcase
        end
    end

`ifdef SIM
    always @(negedge clk) begin
        if (!reset_n) begin
            instr[11:6] <= 0;
            instr[23:18] <= 0;
            instr[31:30] <= 0;
            in1[11:6] <= 0;
            in2[11:6] <= 0;
        end
        else begin
            case (addr)
            0: instr[11: 6] <= io_in;
            1: instr[23:18] <= io_in;
            2: instr[31:30] <= io_in;
            3: in1[11: 6] <= io_in;
            4: in2[11: 6] <= io_in;
            endcase
        end
    end
`else
    generate
        for (i = 0; i < 6; i = i + 1) begin
            sky130_fd_sc_hd__dfrtn_1 instr1ff(.Q(instr[i+6]), .D((addr == 0) ? io_in[i] : instr[i+6]), .CLK_N(clk), .RESET_B(reset_n));
            sky130_fd_sc_hd__dfrtn_1 instr2ff(.Q(instr[i+18]), .D((addr == 1) ? io_in[i] : instr[i+18]), .CLK_N(clk), .RESET_B(reset_n));
            if (i < 2) sky130_fd_sc_hd__dfrtn_1 instr3ff(.Q(instr[i+30]), .D((addr == 2) ? io_in[i] : instr[i+30]), .CLK_N(clk), .RESET_B(reset_n));
            sky130_fd_sc_hd__dfrtn_1 in1ff(.Q(in1[i+6]), .D((addr == 3) ? io_in[i] : in1[i+6]), .CLK_N(clk), .RESET_B(reset_n));
            sky130_fd_sc_hd__dfrtn_1 in2ff(.Q(in2[i+6]), .D((addr == 4) ? io_in[i] : in2[i+6]), .CLK_N(clk), .RESET_B(reset_n));
        end
    endgenerate
`endif

    function [7:0] get_out(input [2:0] addr);
        case (addr)
        2: begin
            get_out[0] = in1_adv;
            get_out[1] = in2_adv;
            get_out[2] = out_valid && !out_select;
            get_out[3] = out_valid && out_select;
            get_out[7:4] = 0;
        end
        4: get_out = pc;
        0: get_out = out[ 7: 0];
        1: get_out = { 4'b0000, out[11: 8] };
        3: get_out = { out[11], seg7_out };
        endcase
    endfunction

    assign io_out = get_out(addr);

endmodule