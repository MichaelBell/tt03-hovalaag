`default_nettype none
`timescale 1ns/1ps

/*
this testbench just instantiates the module and makes some convenient wires
that can be driven / tested by the cocotb test.py
*/

module tb (
    // testbench is controlled by test.py
    input clk,
    input rst,
    input [5:0] data_in,
    output [7:0] data_out
   );

    // this part dumps the trace to a vcd file that can be viewed with GTKWave
    initial begin
        $dumpfile ("tb.vcd");
        $dumpvars (0, tb);
        #1;
    end

    // wire up the inputs and outputs
    wire [7:0] inputs = {data_in[5:0], !rst, clk};
    wire [7:0] outputs;
    assign data_out = outputs;

    // instantiate the DUT
    MichaelBell_hovalaag uut(
`ifdef GL_TEST
        // for gatelevel testing we need to set up the power pins
        .vccd1(1'b1),
        .vssd1(1'b0),
`endif
        .io_in  (inputs),
        .io_out (outputs)
        );

endmodule
