/* Copyright (C) 2023 Michael Bell

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
*/

/* Top module for the Hovalaag Tiny Tapeout
 *
 * IN: 0: CLK
 *     1: RESET_EN
 *   2-7: DATA if RESET_EN false
 *     2: RESET if RESET_EN true
 *     3: RESET address only
 */

module MichaelBell_hovalaag (
  input [7:0] io_in,
  output [7:0] io_out
);
    wire clk = io_in[0];

    wire reset;
    reg reset_rosc;

    reg [3:0] addr;
    reg [3:0] next_addr;

    assign reset = io_in[1] && io_in[2];

    HovalaagWrapper wrapper (
        .clk(clk),
        .reset(reset),
        .reset_rosc(reset_rosc),
        .addr(addr),
        .io_in(io_in[7:2]),
        .io_out(io_out[7:0])
    );

    always @(posedge clk) begin
        if (io_in[1] && io_in[2]) begin
            reset_rosc <= 1'b1;
        end 
        else if (io_in[1] && io_in[4]) begin
            reset_rosc <= 1'b0;
        end

        if (io_in[1] && (io_in[2] || io_in[3])) begin
            next_addr <= 4'h0;
        end
        else begin
            if (next_addr == 9) next_addr <= 0;
            else next_addr <= next_addr + 1;
        end
    end

    always @(negedge clk) begin
        addr <= next_addr;
    end

endmodule